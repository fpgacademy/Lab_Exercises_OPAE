module memory_to_stream_dma_bbb (
		input  wire         clk_clk,                        //              clk.clk
		output wire         csr_waitrequest,                //              csr.waitrequest
		output wire [63:0]  csr_readdata,                   //                 .readdata
		output wire         csr_readdatavalid,              //                 .readdatavalid
		input  wire [0:0]   csr_burstcount,                 //                 .burstcount
		input  wire [63:0]  csr_writedata,                  //                 .writedata
		input  wire [7:0]   csr_address,                    //                 .address
		input  wire         csr_write,                      //                 .write
		input  wire         csr_read,                       //                 .read
		input  wire [7:0]   csr_byteenable,                 //                 .byteenable
		input  wire         csr_debugaccess,                //                 .debugaccess
		input  wire         host_read_waitrequest,          //        host_read.waitrequest
		input  wire [511:0] host_read_readdata,             //                 .readdata
		input  wire         host_read_readdatavalid,        //                 .readdatavalid
		output wire [2:0]   host_read_burstcount,           //                 .burstcount
		output wire [511:0] host_read_writedata,            //                 .writedata
		output wire [47:0]  host_read_address,              //                 .address
		output wire         host_read_write,                //                 .write
		output wire         host_read_read,                 //                 .read
		output wire [63:0]  host_read_byteenable,           //                 .byteenable
		output wire         host_read_debugaccess,          //                 .debugaccess
		output wire [47:0]  descriptor_fetch_address,       // descriptor_fetch.address
		output wire [2:0]   descriptor_fetch_burstcount,    //                 .burstcount
		output wire [63:0]  descriptor_fetch_byteenable,    //                 .byteenable
		output wire         descriptor_fetch_read,          //                 .read
		input  wire [511:0] descriptor_fetch_readdata,      //                 .readdata
		input  wire         descriptor_fetch_readdatavalid, //                 .readdatavalid
		input  wire         descriptor_fetch_waitrequest,   //                 .waitrequest
		output wire [47:0]  descriptor_store_address,       // descriptor_store.address
		output wire [2:0]   descriptor_store_burstcount,    //                 .burstcount
		output wire [63:0]  descriptor_store_byteenable,    //                 .byteenable
		input  wire         descriptor_store_waitrequest,   //                 .waitrequest
		output wire         descriptor_store_write,         //                 .write
		output wire [511:0] descriptor_store_writedata,     //                 .writedata
		input  wire         mem_read_waitrequest,           //         mem_read.waitrequest
		input  wire [511:0] mem_read_readdata,              //                 .readdata
		input  wire         mem_read_readdatavalid,         //                 .readdatavalid
		output wire [2:0]   mem_read_burstcount,            //                 .burstcount
		output wire [511:0] mem_read_writedata,             //                 .writedata
		output wire [47:0]  mem_read_address,               //                 .address
		output wire         mem_read_write,                 //                 .write
		output wire         mem_read_read,                  //                 .read
		output wire [63:0]  mem_read_byteenable,            //                 .byteenable
		output wire         mem_read_debugaccess,           //                 .debugaccess
		output wire [511:0] m2s_st_source_data,             //    m2s_st_source.data
		output wire         m2s_st_source_valid,            //                 .valid
		input  wire         m2s_st_source_ready,            //                 .ready
		output wire         m2s_st_source_startofpacket,    //                 .startofpacket
		output wire         m2s_st_source_endofpacket,      //                 .endofpacket
		output wire [5:0]   m2s_st_source_empty,            //                 .empty
		input  wire         reset_reset                     //            reset.reset
	);
endmodule

